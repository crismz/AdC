//REGFILE

module regfile	(input logic clk,
					 input logic we3,
					 input logic [4:0] ra1,
					 input logic [4:0] ra2,
					 input logic [4:0] wa3,
					 input logic [63:0] wd3,
					 output logic [63:0] rd1,
					 output logic [63:0] rd2);
					 
	logic [63:0] REGS [0:31];
	
	initial 
	begin
		REGS  = '{default:'0};
		for (logic [63-1:0] i = 0; i < 'd31; ++i) REGS[i] = i;
	end
	
	always @(posedge clk)
		if (we3)
			REGS[wa3] <= wd3;

		always_comb begin
			if (we3 && (wa3 != 5'd31)) begin
				if (ra1 == wa3) begin
					rd1 <= wd3;
					rd2 <= (ra2 == 5'd31) ? 64'b0 : REGS[ra2];
				end
				else if (ra2 == wa3) begin
					rd1 <= (ra1 == 5'd31) ? 64'b0 : REGS[ra1];
					rd2 <= wd3;
				end
				else begin
					rd1 <= (ra1 == 5'd31) ? 64'b0 : REGS[ra1];
					rd2 <= (ra2 == 5'd31) ? 64'b0 : REGS[ra2];
				end
			end 
			else begin
				rd1 <= (ra1 == 5'd31) ? 64'b0 : REGS[ra1];
				rd2 <= (ra2 == 5'd31) ? 64'b0 : REGS[ra2];
			end
		end
					 

endmodule